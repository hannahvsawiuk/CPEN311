// Implements a simple Nios II system for the DE-series board.// Inputs:  SW7−0 are parallel port inputs to the Nios II system
//          CLOCK_50 is the system clock
//          KEY[0] is the active-low system reset  // Outputs: LEDR7−0 are parallel port outputs from the Nios II system
module lights (CLOCK_50, SW, KEY, LEDR, HEX0, HEX1);input CLOCK_50; 
input [7:0] SW; 
input [0:0] KEY; 
output [7:0] LEDR;wire [7:0] ledin;output [6:0] HEX0, HEX1;// Instantiate the Nios II system module generated by the Qsys tool: 

nios_system NiosII (   .clk_clk(CLOCK_50),  
   .reset_reset_n(KEY), 
   .switches_export(SW), 
   .leds_export(LEDR),   .ledin_export(ledin));   seven_seg hex0(ledin[3:0], HEX0);seven_seg hex1(ledin[7:4], HEX1);  endmodule